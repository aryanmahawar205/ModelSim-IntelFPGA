//Test Bench for Full Adder

module TB_fullAdder();
wire sum, carry; reg A, B, Cin;

