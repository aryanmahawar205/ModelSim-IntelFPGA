//structural modelling for Full Adder

module exp_str(sum, carry, A, B, Cin);
input A, B, Cin; output sum, carry;
xor g1(sum, A, B, Cin);
wire y1, y2, y3;
and g2(y1, B, Cin);
and g3(y2, A, B);
and g4(y3, A, Cin);
and g5(carry, y1, y2, y3);
endmodule